magic
tech sky130A
timestamp 1723843874
<< metal4 >>
rect 600 500 650 650
rect 850 500 900 650
use sky130_fd_pr__cap_mim_m3_1_BZXSER  sky130_fd_pr__cap_mim_m3_1_BZXSER_0
timestamp 1723843874
transform 1 0 446 0 1 367
box -443 -370 443 370
<< labels >>
flabel metal4 850 500 900 650 0 FreeSans 800 0 0 0 A
port 0 nsew
flabel metal4 600 500 650 650 0 FreeSans 800 0 0 0 B
port 1 nsew
<< end >>
