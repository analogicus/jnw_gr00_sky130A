module JNWG00_CCELL
(
  input wire VDD_1V8,
  inout wire CB,
  inout wire CA,
  input wire CB_1V8,
  input wire CA_1V8,
  input wire VSS,
);

endmodule
