*Model comparator
.subckt JNWG00_CMP SWAP_1V8 VN VP VSS ZERO_1V8 PWRUP_1V8 CMPO VDD_1V8 IBN

I1 0 VCN 5u
x1 VCN VCN VSS VSS JNWATR_NCH_2C1F2
x2 IBN VCN VSS VSS JNWATR_NCH_2C1F2
C1 VP 0 100f
C2 VN 0 100f
E1 CMPO VSS value={v(VDD_1V8)*(tanh(10000*(v(vp)-v(vn)))+1)/2) }
.ends
