module JNWG00_CCELL
(
  input wire VDD_1V8,
  inout wire CA,
  input wire CA_1V8,
  input wire VSS,
  inout wire CB,
  input wire CB_1V8
);

endmodule
