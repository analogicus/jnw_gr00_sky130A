magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 0 0
use JNWATR_PCH_8C5F0 x11[2:0] ../JNW_ATR_SKY130A
transform 1 0 0 0 1 0
box 0 0 0 0
use JNWATR_PCH_8C5F0 x11[2:0] ../JNW_ATR_SKY130A
transform 1 0 0 0 1 400
box 0 400 0 400
use JNWATR_PCH_8C5F0 x14[2:0] ../JNW_ATR_SKY130A
transform 1 0 704 0 1 0
box 704 0 704 0
use JNWATR_PCH_8C5F0 x14[2:0] ../JNW_ATR_SKY130A
transform 1 0 704 0 1 400
box 704 400 704 400
use JNWATR_PCH_8C1F2 x15[2:0] ../JNW_ATR_SKY130A
transform 1 0 1408 0 1 0
box 1408 0 1408 0
use JNWATR_PCH_8C1F2 x15[2:0] ../JNW_ATR_SKY130A
transform 1 0 1408 0 1 400
box 1408 400 1408 400
use JNWATR_PCH_8C1F2 x16[2:0] ../JNW_ATR_SKY130A
transform 1 0 2112 0 1 0
box 2112 0 2112 0
use JNWATR_PCH_8C1F2 x16[2:0] ../JNW_ATR_SKY130A
transform 1 0 2112 0 1 400
box 2112 400 2112 400
use JNWATR_NCH_2C1F2 x17[3:0] ../JNW_ATR_SKY130A
transform 1 0 2816 0 1 0
box 2816 0 2816 0
use JNWATR_NCH_2C1F2 x17[3:0] ../JNW_ATR_SKY130A
transform 1 0 2816 0 1 400
box 2816 400 2816 400
use JNWATR_NCH_2C1F2 x17[3:0] ../JNW_ATR_SKY130A
transform 1 0 2816 0 1 800
box 2816 800 2816 800
use JNWATR_NCH_2C5F0 x18[3:0] ../JNW_ATR_SKY130A
transform 1 0 3328 0 1 0
box 3328 0 3328 0
use JNWATR_NCH_2C5F0 x18[3:0] ../JNW_ATR_SKY130A
transform 1 0 3328 0 1 400
box 3328 400 3328 400
use JNWATR_NCH_2C5F0 x18[3:0] ../JNW_ATR_SKY130A
transform 1 0 3328 0 1 800
box 3328 800 3328 800
use JNWATR_NCH_2C1F2 x19[3:0] ../JNW_ATR_SKY130A
transform 1 0 3840 0 1 0
box 3840 0 3840 0
use JNWATR_NCH_2C1F2 x19[3:0] ../JNW_ATR_SKY130A
transform 1 0 3840 0 1 400
box 3840 400 3840 400
use JNWATR_NCH_2C1F2 x19[3:0] ../JNW_ATR_SKY130A
transform 1 0 3840 0 1 800
box 3840 800 3840 800
use JNWATR_NCH_2C5F0 x20[3:0] ../JNW_ATR_SKY130A
transform 1 0 4352 0 1 0
box 4352 0 4352 0
use JNWATR_NCH_2C5F0 x20[3:0] ../JNW_ATR_SKY130A
transform 1 0 4352 0 1 400
box 4352 400 4352 400
use JNWATR_NCH_2C5F0 x20[3:0] ../JNW_ATR_SKY130A
transform 1 0 4352 0 1 800
box 4352 800 4352 800
use JNWATR_NCH_2C5F0 x22 ../JNW_ATR_SKY130A
transform 1 0 4864 0 1 0
box 4864 0 4864 0
use JNWATR_PCH_8C5F0 x23 ../JNW_ATR_SKY130A
transform 1 0 5376 0 1 0
box 5376 0 5376 0
use JNWATR_PCH_8C1F2 x24 ../JNW_ATR_SKY130A
transform 1 0 6080 0 1 0
box 6080 0 6080 0
use JNWATR_NCH_2C1F2 x25 ../JNW_ATR_SKY130A
transform 1 0 6784 0 1 0
box 6784 0 6784 0
use JNWTR_RPPO16 x26 ../JNW_TR_SKY130A
transform 1 0 7296 0 1 0
box 7296 0 7296 0
use JNWTR_RPPO16 x27 ../JNW_TR_SKY130A
transform 1 0 9532 0 1 0
box 9532 0 9532 0
use JNWATR_NCH_2C5F0 x28 ../JNW_ATR_SKY130A
transform 1 0 11768 0 1 0
box 11768 0 11768 0
use JNWATR_NCH_2C1F2 x29 ../JNW_ATR_SKY130A
transform 1 0 12280 0 1 0
box 12280 0 12280 0
use JNWATR_PCH_4C1F2 x30 ../JNW_ATR_SKY130A
transform 1 0 12792 0 1 0
box 12792 0 12792 0
use JNWTR_RPPO4 x31 ../JNW_TR_SKY130A
transform 1 0 13368 0 1 0
box 13368 0 13368 0
use JNWATR_PCH_8C1F2 x32 ../JNW_ATR_SKY130A
transform 1 0 14308 0 1 0
box 14308 0 14308 0
use JNWATR_NCH_2C1F2 x33 ../JNW_ATR_SKY130A
transform 1 0 15012 0 1 0
box 15012 0 15012 0
use JNWTR_IVX1_CV x34 ../JNW_TR_SKY130A
transform 1 0 15524 0 1 0
box 15524 0 15524 0
use JNWTR_RPPO8 x11 ../JNW_TR_SKY130A
transform 1 0 16514 0 1 0
box 16514 0 16514 0
use JNWATR_PCH_8C5F0 x35 ../JNW_ATR_SKY130A
transform 1 0 17886 0 1 0
box 17886 0 17886 0
use JNWATR_NCH_2C5F0 x36 ../JNW_ATR_SKY130A
transform 1 0 18590 0 1 0
box 18590 0 18590 0
use JNWATR_PCH_12C1F2 x3[3:0] ../JNW_ATR_SKY130A
transform 1 0 19102 0 1 0
box 19102 0 19102 0
use JNWATR_PCH_12C1F2 x3[3:0] ../JNW_ATR_SKY130A
transform 1 0 19102 0 1 400
box 19102 400 19102 400
use JNWATR_PCH_12C1F2 x3[3:0] ../JNW_ATR_SKY130A
transform 1 0 19102 0 1 800
box 19102 800 19102 800
use JNWATR_PCH_12C1F2 x4[3:0] ../JNW_ATR_SKY130A
transform 1 0 19934 0 1 0
box 19934 0 19934 0
use JNWATR_PCH_12C1F2 x4[3:0] ../JNW_ATR_SKY130A
transform 1 0 19934 0 1 400
box 19934 400 19934 400
use JNWATR_PCH_12C1F2 x4[3:0] ../JNW_ATR_SKY130A
transform 1 0 19934 0 1 800
box 19934 800 19934 800
use JNWATR_PCH_8C5F0 x1[1:0] ../JNW_ATR_SKY130A
transform 1 0 20766 0 1 0
box 20766 0 20766 0
use JNWATR_NCH_2C5F0 x1 ../JNW_ATR_SKY130A
transform 1 0 21470 0 1 0
box 21470 0 21470 0
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130A
transform 1 0 21982 0 1 0
box 21982 0 21982 0
use JNWTR_RPPO16 x6 ../JNW_TR_SKY130A
transform 1 0 22494 0 1 0
box 22494 0 22494 0
use JNWTR_RPPO16 x7 ../JNW_TR_SKY130A
transform 1 0 24730 0 1 0
box 24730 0 24730 0
use JNWATR_NCH_2C1F2 x8 ../JNW_ATR_SKY130A
transform 1 0 26966 0 1 0
box 26966 0 26966 0
use JNWATR_NCH_2C1F2 x18 ../JNW_ATR_SKY130A
transform 1 0 27478 0 1 0
box 27478 0 27478 0
use JNWTR_IVX1_CV x38 ../JNW_TR_SKY130A
transform 1 0 27990 0 1 0
box 27990 0 27990 0
use JNWATR_PCH_2C1F2 x4 ../JNW_ATR_SKY130A
transform 1 0 28980 0 1 0
box 28980 0 28980 0
use JNWATR_PCH_2C1F2 x5 ../JNW_ATR_SKY130A
transform 1 0 29492 0 1 0
box 29492 0 29492 0
use JNWATR_PCH_2C5F0 x3 ../JNW_ATR_SKY130A
transform 1 0 30004 0 1 0
box 30004 0 30004 0
use JNWTR_RPPO8 x39 ../JNW_TR_SKY130A
transform 1 0 30516 0 1 0
box 30516 0 30516 0
use JNWTR_IVX1_CV x40 ../JNW_TR_SKY130A
transform 1 0 31888 0 1 0
box 31888 0 31888 0
use JNWTR_IVX1_CV x16 ../JNW_TR_SKY130A
transform 1 0 32878 0 1 0
box 32878 0 32878 0
use JNWTR_IVX1_CV x14 ../JNW_TR_SKY130A
transform 1 0 33868 0 1 0
box 33868 0 33868 0
use JNWTR_IVX1_CV x41 ../JNW_TR_SKY130A
transform 1 0 34858 0 1 0
box 34858 0 34858 0
use JNWTR_IVX1_CV x42 ../JNW_TR_SKY130A
transform 1 0 35848 0 1 0
box 35848 0 35848 0
use JNWTR_IVX1_CV x17 ../JNW_TR_SKY130A
transform 1 0 36838 0 1 0
box 36838 0 36838 0
use JNWTR_IVX1_CV x19 ../JNW_TR_SKY130A
transform 1 0 37828 0 1 0
box 37828 0 37828 0
use JNWTR_IVX1_CV x20 ../JNW_TR_SKY130A
transform 1 0 38818 0 1 0
box 38818 0 38818 0
use JNWTR_IVX1_CV x21 ../JNW_TR_SKY130A
transform 1 0 39808 0 1 0
box 39808 0 39808 0
use JNWTR_NCHDL x12[1:0] ../JNW_TR_SKY130A
transform 1 0 40798 0 1 0
box 40798 0 40798 0
use JNWTR_NCHDL x2[1:0] ../JNW_TR_SKY130A
transform 1 0 41293 0 1 0
box 41293 0 41293 0
use JNWTR_NCHDL x12 ../JNW_TR_SKY130A
transform 1 0 41788 0 1 0
box 41788 0 41788 0
use JNWTR_NCHDL x13 ../JNW_TR_SKY130A
transform 1 0 42283 0 1 0
box 42283 0 42283 0
use JNWTR_CAPX1 x37[1:0] ../JNW_TR_SKY130A
transform 1 0 42778 0 1 0
box 42778 0 42778 0
use JNWTR_CAPX1 x6[1:0] ../JNW_TR_SKY130A
transform 1 0 43318 0 1 0
box 43318 0 43318 0
use JNWTR_CAPX1 x7[1:0] ../JNW_TR_SKY130A
transform 1 0 43858 0 1 0
box 43858 0 43858 0
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 0
box 44398 0 44398 0
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 540
box 44398 540 44398 540
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 1080
box 44398 1080 44398 1080
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 1620
box 44398 1620 44398 1620
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 2160
box 44398 2160 44398 2160
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 2700
box 44398 2700 44398 2700
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 3240
box 44398 3240 44398 3240
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 3780
box 44398 3780 44398 3780
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 4320
box 44398 4320 44398 4320
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 4860
box 44398 4860 44398 4860
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 5400
box 44398 5400 44398 5400
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 5940
box 44398 5940 44398 5940
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 6480
box 44398 6480 44398 6480
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 7020
box 44398 7020 44398 7020
use JNWTR_CAPX1 x5[15:0] ../JNW_TR_SKY130A
transform 1 0 44398 0 1 7560
box 44398 7560 44398 7560
use JNWTR_TGX2_CV x10 ../JNW_TR_SKY130A
transform 1 0 44938 0 1 0
box 44938 0 44938 0
use JNWTR_TGX2_CV x9 ../JNW_TR_SKY130A
transform 1 0 45928 0 1 0
box 45928 0 45928 0
<< labels >>
<< properties >>
<< end >>
