module JNWG00_CMP
(
 input wire  VDD_1V8,
 input wire  VSS,
 input wire  VP,
 output wire CMPO,
 input wire  VN,
 input wire  SWAP_1V8,
 input wire  PWRUP_1V8,
 input wire  ZERO_1V8
);


endmodule
