magic
tech sky130A
magscale 1 1
timestamp 1723759200
<< checkpaint >>
rect 0 0 0 0
use JNWATR_PCH_8C5F0 x11[2:0] ../JNW_ATR_SKY130NM
transform 1 0 0 0 1 0
box 0 0 0 0
use JNWATR_PCH_8C5F0 x11[2:0] ../JNW_ATR_SKY130NM
transform 1 0 0 0 1 400
box 0 400 0 400
use JNWATR_PCH_8C5F0 x14[2:0] ../JNW_ATR_SKY130NM
transform 1 0 704 0 1 0
box 704 0 704 0
use JNWATR_PCH_8C5F0 x14[2:0] ../JNW_ATR_SKY130NM
transform 1 0 704 0 1 400
box 704 400 704 400
use JNWATR_PCH_8C1F2 x15[2:0] ../JNW_ATR_SKY130NM
transform 1 0 1408 0 1 0
box 1408 0 1408 0
use JNWATR_PCH_8C1F2 x15[2:0] ../JNW_ATR_SKY130NM
transform 1 0 1408 0 1 400
box 1408 400 1408 400
use JNWATR_PCH_8C1F2 x16[2:0] ../JNW_ATR_SKY130NM
transform 1 0 2112 0 1 0
box 2112 0 2112 0
use JNWATR_PCH_8C1F2 x16[2:0] ../JNW_ATR_SKY130NM
transform 1 0 2112 0 1 400
box 2112 400 2112 400
use JNWATR_NCH_2C1F2 x17[3:0] ../JNW_ATR_SKY130NM
transform 1 0 2816 0 1 0
box 2816 0 2816 0
use JNWATR_NCH_2C1F2 x17[3:0] ../JNW_ATR_SKY130NM
transform 1 0 2816 0 1 400
box 2816 400 2816 400
use JNWATR_NCH_2C1F2 x17[3:0] ../JNW_ATR_SKY130NM
transform 1 0 2816 0 1 800
box 2816 800 2816 800
use JNWATR_NCH_2C5F0 x18[3:0] ../JNW_ATR_SKY130NM
transform 1 0 3328 0 1 0
box 3328 0 3328 0
use JNWATR_NCH_2C5F0 x18[3:0] ../JNW_ATR_SKY130NM
transform 1 0 3328 0 1 400
box 3328 400 3328 400
use JNWATR_NCH_2C5F0 x18[3:0] ../JNW_ATR_SKY130NM
transform 1 0 3328 0 1 800
box 3328 800 3328 800
use JNWATR_NCH_2C1F2 x19[3:0] ../JNW_ATR_SKY130NM
transform 1 0 3840 0 1 0
box 3840 0 3840 0
use JNWATR_NCH_2C1F2 x19[3:0] ../JNW_ATR_SKY130NM
transform 1 0 3840 0 1 400
box 3840 400 3840 400
use JNWATR_NCH_2C1F2 x19[3:0] ../JNW_ATR_SKY130NM
transform 1 0 3840 0 1 800
box 3840 800 3840 800
use JNWATR_NCH_2C5F0 x20[3:0] ../JNW_ATR_SKY130NM
transform 1 0 4352 0 1 0
box 4352 0 4352 0
use JNWATR_NCH_2C5F0 x20[3:0] ../JNW_ATR_SKY130NM
transform 1 0 4352 0 1 400
box 4352 400 4352 400
use JNWATR_NCH_2C5F0 x20[3:0] ../JNW_ATR_SKY130NM
transform 1 0 4352 0 1 800
box 4352 800 4352 800
use JNWATR_NCH_2C5F0 x22 ../JNW_ATR_SKY130NM
transform 1 0 4864 0 1 0
box 4864 0 4864 0
use JNWATR_PCH_8C5F0 x23 ../JNW_ATR_SKY130NM
transform 1 0 5376 0 1 0
box 5376 0 5376 0
use JNWATR_PCH_8C1F2 x24 ../JNW_ATR_SKY130NM
transform 1 0 6080 0 1 0
box 6080 0 6080 0
use JNWATR_NCH_2C1F2 x25 ../JNW_ATR_SKY130NM
transform 1 0 6784 0 1 0
box 6784 0 6784 0
use SUNTR_RPPO16 x26 ../SUN_TR_SKY130NM
transform 1 0 7296 0 1 0
box 7296 0 7296 0
use SUNTR_RPPO16 x27 ../SUN_TR_SKY130NM
transform 1 0 11656 0 1 0
box 11656 0 11656 0
use JNWATR_NCH_2C5F0 x28 ../JNW_ATR_SKY130NM
transform 1 0 16016 0 1 0
box 16016 0 16016 0
use JNWATR_NCH_2C1F2 x29 ../JNW_ATR_SKY130NM
transform 1 0 16528 0 1 0
box 16528 0 16528 0
use JNWATR_PCH_4C1F2 x30 ../JNW_ATR_SKY130NM
transform 1 0 17040 0 1 0
box 17040 0 17040 0
use SUNTR_RPPO4 x31 ../SUN_TR_SKY130NM
transform 1 0 17616 0 1 0
box 17616 0 17616 0
use JNWATR_PCH_8C1F2 x32 ../JNW_ATR_SKY130NM
transform 1 0 19384 0 1 0
box 19384 0 19384 0
use JNWATR_NCH_2C1F2 x33 ../JNW_ATR_SKY130NM
transform 1 0 20088 0 1 0
box 20088 0 20088 0
use SUNTR_IVX1_CV x34 ../SUN_TR_SKY130NM
transform 1 0 20600 0 1 0
box 20600 0 20600 0
use SUNTR_RPPO8 x11 ../SUN_TR_SKY130NM
transform 1 0 21860 0 1 0
box 21860 0 21860 0
use JNWATR_PCH_8C5F0 x35 ../JNW_ATR_SKY130NM
transform 1 0 24492 0 1 0
box 24492 0 24492 0
use JNWATR_NCH_2C5F0 x36 ../JNW_ATR_SKY130NM
transform 1 0 25196 0 1 0
box 25196 0 25196 0
use JNWATR_PCH_12C1F2 x3[3:0] ../JNW_ATR_SKY130NM
transform 1 0 25708 0 1 0
box 25708 0 25708 0
use JNWATR_PCH_12C1F2 x3[3:0] ../JNW_ATR_SKY130NM
transform 1 0 25708 0 1 400
box 25708 400 25708 400
use JNWATR_PCH_12C1F2 x3[3:0] ../JNW_ATR_SKY130NM
transform 1 0 25708 0 1 800
box 25708 800 25708 800
use JNWATR_PCH_12C1F2 x4[3:0] ../JNW_ATR_SKY130NM
transform 1 0 26540 0 1 0
box 26540 0 26540 0
use JNWATR_PCH_12C1F2 x4[3:0] ../JNW_ATR_SKY130NM
transform 1 0 26540 0 1 400
box 26540 400 26540 400
use JNWATR_PCH_12C1F2 x4[3:0] ../JNW_ATR_SKY130NM
transform 1 0 26540 0 1 800
box 26540 800 26540 800
use JNWATR_PCH_8C5F0 x1[1:0] ../JNW_ATR_SKY130NM
transform 1 0 27372 0 1 0
box 27372 0 27372 0
use JNWATR_NCH_2C5F0 x1 ../JNW_ATR_SKY130NM
transform 1 0 28076 0 1 0
box 28076 0 28076 0
use JNWATR_NCH_2C1F2 x2 ../JNW_ATR_SKY130NM
transform 1 0 28588 0 1 0
box 28588 0 28588 0
use SUNTR_RPPO16 x6 ../SUN_TR_SKY130NM
transform 1 0 29100 0 1 0
box 29100 0 29100 0
use SUNTR_RPPO16 x7 ../SUN_TR_SKY130NM
transform 1 0 33460 0 1 0
box 33460 0 33460 0
use JNWATR_NCH_2C1F2 x8 ../JNW_ATR_SKY130NM
transform 1 0 37820 0 1 0
box 37820 0 37820 0
use JNWATR_NCH_2C1F2 x18 ../JNW_ATR_SKY130NM
transform 1 0 38332 0 1 0
box 38332 0 38332 0
use SUNTR_IVX1_CV x38 ../SUN_TR_SKY130NM
transform 1 0 38844 0 1 0
box 38844 0 38844 0
use JNWATR_PCH_2C1F2 x4 ../JNW_ATR_SKY130NM
transform 1 0 40104 0 1 0
box 40104 0 40104 0
use JNWATR_PCH_2C1F2 x5 ../JNW_ATR_SKY130NM
transform 1 0 40616 0 1 0
box 40616 0 40616 0
use JNWATR_PCH_2C5F0 x3 ../JNW_ATR_SKY130NM
transform 1 0 41128 0 1 0
box 41128 0 41128 0
use SUNTR_RPPO8 x39 ../SUN_TR_SKY130NM
transform 1 0 41640 0 1 0
box 41640 0 41640 0
use SUNTR_IVX1_CV x40 ../SUN_TR_SKY130NM
transform 1 0 44272 0 1 0
box 44272 0 44272 0
use JNWG00_TG x10 ../JNW_GR00_SKY130NM
transform 1 0 45532 0 1 0
box 45532 0 45532 0
use SUNTR_IVX1_CV x16 ../SUN_TR_SKY130NM
transform 1 0 45532 0 1 0
box 45532 0 45532 0
use SUNTR_IVX1_CV x14 ../SUN_TR_SKY130NM
transform 1 0 46792 0 1 0
box 46792 0 46792 0
use SUNTR_IVX1_CV x41 ../SUN_TR_SKY130NM
transform 1 0 48052 0 1 0
box 48052 0 48052 0
use SUNTR_IVX1_CV x42 ../SUN_TR_SKY130NM
transform 1 0 49312 0 1 0
box 49312 0 49312 0
use JNWG00_TG x9 ../JNW_GR00_SKY130NM
transform 1 0 50572 0 1 0
box 50572 0 50572 0
use SUNTR_IVX1_CV x17 ../SUN_TR_SKY130NM
transform 1 0 50572 0 1 0
box 50572 0 50572 0
use SUNTR_IVX1_CV x19 ../SUN_TR_SKY130NM
transform 1 0 51832 0 1 0
box 51832 0 51832 0
use SUNTR_IVX1_CV x20 ../SUN_TR_SKY130NM
transform 1 0 53092 0 1 0
box 53092 0 53092 0
use SUNTR_IVX1_CV x21 ../SUN_TR_SKY130NM
transform 1 0 54352 0 1 0
box 54352 0 54352 0
use SUNTR_NCHDL x12[1:0] ../SUN_TR_SKY130NM
transform 1 0 55612 0 1 0
box 55612 0 55612 0
use SUNTR_NCHDL x2[1:0] ../SUN_TR_SKY130NM
transform 1 0 56242 0 1 0
box 56242 0 56242 0
use SUNTR_NCHDL x12 ../SUN_TR_SKY130NM
transform 1 0 56872 0 1 0
box 56872 0 56872 0
use SUNTR_NCHDL x13 ../SUN_TR_SKY130NM
transform 1 0 57502 0 1 0
box 57502 0 57502 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x5[9:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x15 ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x37[1:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
use JNWG00_UCAP x43[1:0] ../JNW_GR00_SKY130NM
transform 1 0 58132 0 1 0
box 58132 0 58132 0
<< labels >>
<< properties >>
<< end >>
