module JNWG00_IDAC
(
  input wire [7:0] IBF,
  input wire [7:0] IB,
  input wire VDD_1V8,
  inout wire [3:0] IDAC_O,
  input wire [3:0] IBO_N_1V8,
  input wire PWRUP_1V8,
  input wire VSS
);

   endmodule
