module JNWG00_BDAC
(
  input wire [7:0] BD_1V8,
  inout wire VD,
  input wire VSS,
  input wire RES_N_1V8,
  input wire R_IBPS_1V8
);

endmodule // JNWG00_BDAC
